module EXP6 (

input clk, // Clock input

input reset, // Reset input (active high)

output [3:0] q // 4-bit output

);

// Internal signals for flip-flops

reg [3:0] q_int;

// Assign internal register to output

assign q = q_int;

always @(posedge clk or posedge reset) begin

if (reset)

q_int[0] <= 1'b0; // Reset the first bit to 0

else

q_int[0] <= ~q_int[0]; // Toggle the first bit on clock edge

end

// Generate the other flip-flops based on the output of the previous one

genvar i;

generate

for (i = 1; i < 4; i = i + 1) begin : ripple

always @(posedge q_int[i-1] or posedge reset) begin

if (reset)

q_int[i] <= 1'b0; // Reset the bit to 0

else

q_int[i] <= ~q_int[i]; // Toggle the bit on clock edge of previous stage

end

end

endgenerate

endmodule